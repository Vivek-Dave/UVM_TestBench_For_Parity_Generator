
interface intf();
    // ------------------- port declaration-------------------------------------
    logic  [7:0] data;
    logic even_parity;
    logic  odd_parity;
    //--------------------------------------------------------------------------        
endinterface

